module round_robin #(
    parameter NUM_REQUEST = 4
)(
    input logic clk,
    input logic rst_n,
    // input
    
);
    
endmodule